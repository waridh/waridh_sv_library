module microaddr_counter(
  input logic clk,
  input logic reset,
  input microaddr::cmd cmd,
  input logic[10:0] load_addr,
  output logic[10:0] addr
);


endmodule
